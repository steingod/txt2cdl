netcdf template_bio {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 
// $Id: template_bio.cdl,v 1.6 2010-06-03 22:10:41 steingod Exp $

dimensions:
    depth = +ndepths; 
    stations = +nstations;
    str25 = 25;

variables:
    char stid(stations,str25);
    	stid:long_name = "Station identifier";
    double time(stations);
	time:long_name = "time in UTC the station was taken";
	time:short_name = "time";
	time:standard_name = "time";
	time:units = "seconds since 1970-01-01 00:00:00 UTC";
	time:axis = "T";
    float latitude(stations);
	latitude:long_name = "geographical latitude in degrees North";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.;
	latitude:valid_max = 90.;
    float longitude(stations);
	longitude:long_name = "geographical longitude in degrees East";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.;
	longitude:valid_max = 180.;
    float depth(depth);
	depth:long_name = "Depth below sea surface in meter";
	depth:short_name = "depth";
	depth:standard_name = "depth";
	depth:units = "m";
	depth:valid_min = 0.;
	depth:valid_max = 15000.;
	depth:positive = "down";
	depth:axis = "Y";
    float no3no2(stations,depth);
	no3no2:standard_name = "mole_concentration_of_ phosphate_in_sea_water";
	no3no2:long_name = "Nitrate plus nitrite concentration";
	no3no2:short_name = "no3no2";
	no3no2:_FillValue = 9999.f;
	no3no2:units = "micromol L-1";
	no3no2:coordinates = "time longitude latitude depth";
    float no3no2_stdev(stations,depth);
	no3no2_stdev:long_name = "Phospate concentration standard deviation";
	no3no2_stdev:short_name = "no3no2_stdev";
	no3no2_stdev:_FillValue = 9999.f;
	no3no2_stdev:units = "micromol L-1";
	no3no2_stdev:coordinates = "time longitude latitude depth";
    float PO4(stations,depth);
	PO4:standard_name = "mole_concentration_of_ phosphate_in_sea_water";
	PO4:long_name = "Phosphate concentration";
	PO4:short_name = "PO4";
	PO4:_FillValue = 9999.f;
	PO4:units = "micromol L-1";
	PO4:coordinates = "time longitude latitude depth";
    float PO4_stdev(stations,depth);
	PO4_stdev:long_name = "Phospate concentration standard deviation";
	PO4_stdev:short_name = "PO4_stdev";
	PO4_stdev:_FillValue = 9999.f;
	PO4_stdev:units = "micromol L-1";
	PO4_stdev:coordinates = "time longitude latitude depth";
    float sioh4(stations,depth);
	sioh4:standard_name = "mole_concentration_of_silicate_in_sea_water";
	sioh4:long_name = "Silicate concentration";
	sioh4:short_name = "sioh4";
	sioh4:_FillValue = 9999.f;
	sioh4:units = "micromol L-1";
	sioh4:coordinates = "time longitude latitude depth";
    float sioh4_stdev(stations,depth);
	sioh4_stdev:long_name = "Silicate concentration standard deviation";
	sioh4_stdev:short_name = "sioh4_stdev";
	sioh4_stdev:_FillValue = 9999.f;
	sioh4_stdev:units = "micromol L-1";
	sioh4_stdev:coordinates = "time longitude latitude depth";
    float chl-a(stations,depth);
	chl-a:long_name = "Chlorophyll-A";
	chl-a:short_name = "chl-a";
	chl-a:_FillValue = 9999.f;
	chl-a:units = "milligram liter-1";
	chl-a:coordinates = "time longitude latitude depth";
    float chl-a_stdev(stations,depth);
	chl-a_stdev:long_name = "Chlorophyll-A standard deviation";
	chl-a_stdev:short_name = "chl-a stdev";
	chl-a_stdev:_FillValue = 9999.f;
	chl-a_stdev:units = "milligram m-2 day-2";
	chl-a_stdev:coordinates = "time longitude latitude depth";
    float phaeopigment(stations,depth);
	phaeopigment:long_name = "Phaeopigment";
	phaeopigment:short_name = "phaeopigment";
	phaeopigment:_FillValue = 9999.f;
	phaeopigment:units = "milligram liter-1";
	phaeopigment:coordinates = "time longitude latitude depth";
    float phaeopigment_stdev(stations,depth);
	phaeopigment_stdev:long_name = "Phaeopigment standard deviation";
	phaeopigment_stdev:short_name = "phaeopigment stdev";
	phaeopigment_stdev:_FillValue = 9999.f;
	phaeopigment_stdev:units = "milligram liter-1";
	phaeopigment_stdev:coordinates = "time longitude latitude depth";
    float POC(stations,depth);
	POC:long_name = "Particulate Organic Carbon";
	POC:short_name = "POC";
	POC:_FillValue = 9999.f;
	POC:units = "milligram liter-1";
	POC:coordinates = "time longitude latitude depth";
    float POC_stdev(stations,depth);
	POC_stdev:long_name = "Particulate Organic Carbon standard deviation";
	POC_stdev:short_name = "POC_stdev";
	POC_stdev:_FillValue = 9999.f;
	POC_stdev:units = "milligram liter-1";
	POC_stdev:coordinates = "time longitude latitude depth";
    float PON(stations,depth);
	PON:long_name = "Particulate Organic Nitrogen";
	PON:short_name = "PON";
	PON:_FillValue = 9999.f;
	PON:units = "milligram liter-1";
	PON:coordinates = "time longitude latitude depth";
    float PON_stdev(stations,depth);
	PON_stdev:long_name = "Particulate Organic Nitrogen standard deviation";
	PON_stdev:short_name = "PON_stdev";
	PON_stdev:_FillValue = 9999.f;
	PON_stdev:units = "milligram liter-1";
	PON_stdev:coordinates = "time longitude latitude depth";

// global attributes
	:Conventions = "CF-1.4";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; 
	:topiccategory = "+topic"; 
	:keywords = "+keyw"; 
	:gcmd_keywords = "+gcmdkeyw"; 
	:area = "+area"; 
	:activity_type = "+activity_type";
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:product_name = "+pname";
	:Platform_name = "+vessel";
	:project_name = "+project_name";
	:start_date = "+start_date";
	:stop_date = "+stop_date";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +slat;
	:northernmost_latitude = +nlat;
	:westernmost_longitude = +wlon;
	:easternmost_longitude = +elon;
	:quality_statement = "+qual";

data:
    stid = +stid;
    time =  +time;
    latitude = +lat;
    longitude = +lon;
    depth = +depth;
    no3no2 = +no3no2;
    no3no2_stdev = +no3no2_stdev;
    PO4 = +po4;
    PO4_stdev = +po4_stdev;
    sioh4 = +sioh4;
    sioh4_stdev = +sioh4_stdev;
    chl-a = +chl-a;
    chl-a_stdev = +chl-a_stdev;
    phaeopigment = +pigm;
    phaeopigment_stdev = +pigm_stdev;
    POC = +poc;
    POC_stdev = +poc_stdev;
    PON = +pon;
    PON_stdev = +pon_stdev;
}
