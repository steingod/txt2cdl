netcdf template_bio {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 
// $Id: template_biomassmeso.cdl,v 1.1 2011-01-17 20:43:12 steingod Exp $

dimensions:
    depth = +ndepths; 
    stations = +nstations;
    str25 = 25;

variables:
    char stid(stations,str25);
    	stid:long_name = "Station_identifier";
    double time(stations);
	time:long_name = "time_in_UTC_the_station_was_taken";
	time:short_name = "time";
	time:standard_name = "time";
	time:units = "seconds since 1970-01-01 00:00:00 UTC";
	time:axis = "T";
    float latitude(stations);
	latitude:long_name = "geographical_latitude_in_degrees_North";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.;
	latitude:valid_max = 90.;
    float longitude(stations);
	longitude:long_name = "geographical_longitude_in_degrees_East";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.;
	longitude:valid_max = 180.;
    float depth(depth);
	depth:long_name = "Depth_below_sea_surface_in_meter";
	depth:short_name = "depth";
	depth:standard_name = "depth";
	depth:units = "m";
	depth:valid_min = 0.;
	depth:valid_max = 15000.;
	depth:positive = "down";
	depth:axis = "Y";
    float biomass(stations,depth);
	//biomass:standard_name = "";
	biomass:long_name = "integrated_mesozooplankton_biomass_expressed_as_Carbon";
	biomass:short_name = "biomass";
	biomass:_FillValue = 9999.f;
	biomass:units = "microgram meter-2";
	biomass:coordinates = "time longitude latitude depth";

// global attributes
	:Conventions = "CF-1.4";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; 
	:topiccategory = "+topic"; 
	:keywords = "+keyw"; 
	:gcmd_keywords = "+gcmdkeyw"; 
	:area = "+area"; 
	:activity_type = "+activity";
	:operational_status = "+opstatus";
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:product_name = "+pname";
	:Platform_name = "+vessel";
	:project_name = "+project_name";
	:start_date = "+start_date";
	:stop_date = "+stop_date";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +slat;
	:northernmost_latitude = +nlat;
	:westernmost_longitude = +wlon;
	:easternmost_longitude = +elon;
	:quality_statement = "+qual";

data:
    stid = +stid;
    time =  +time;
    latitude = +lat;
    longitude = +lon;
    depth = +depth;
    biomass = +biomass;
}
