netcdf template_ctd {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 
// $Id: template_ctd_oxygen.cdl,v 1.1 2009-10-06 15:33:48 steingod Exp $

dimensions:
    time = unlimited; //
    n_levels = +nvalues; // maximum number of levels (depth)
    stations = 1;

variables:
    double time(time);
	time:long_name = "time" ;
	time:short_name = "time" ;
	time:standard_name = "time" ;
	time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
	time:axis = "T";
    float latitude(stations);
	latitude:long_name = "latitude";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.;
	latitude:valid_max = 90.;
    float longitude(stations);
	longitude:long_name = "longitude";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.;
	longitude:valid_max = 180.;
    float pres(n_levels);
	pres:long_name = "Sea Water Pressure";
	pres:short_name = "Pressure";
	pres:standard_name = "sea_water_pressure";
	pres:units = "dbar";
	pres:valid_min = 0.;
	pres:valid_max = 15000.;
    float temp(n_levels);
	temp:long_name = "Ocean temperature (ITS-90 deg. C)";
	temp:short_name = "temperature";
	temp:_FillValue = 9999.f;
	temp:units = "degrees Celsius";
    float cond(n_levels);
	cond:long_name = "Ocean conductivity (S/m)";
	cond:short_name = "conductivity";
	cond:standard_name = "sea_water_electrical_conductivity";
	cond:_FillValue = 9999.f;
	cond:units = "S/m";
    float psal(n_levels);
	psal:long_name = "Practical salinity (PSU/sal00)";
	psal:short_name = "salinity";
	psal:standard_name = "sea_water_salinity";
	psal:_FillValue = 9999.f;
	psal:units = "";
    float o2(n_levels);
	o2:long_name = "oxygen content";
	o2:short_name = "oxygen";
	o2:standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water";
	o2:_FillValue = 9999.f;
	o2:units = "micromol kg-1";
	o2:axis = "x";

// global attributes
	:Conventions = "CF-1.0";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; // Add text if wanted
	:topiccategory = "+topic"; // Blank separated list
	:keywords = "+keyw"; // Blank separated list
	:gcmd_keywords = "+gcmdkeyw"; // Newline separated list
	:area = "+area"; // Comma separated list, see http://damocles.met.no/
	:activity_type = "+activity_type";
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:product_name = "+pname";
	:Platform_name = "+vessel";
	:project_name = "+project_name";
	:start_date = "+start_date";
	:stop_date = "+stop_date";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +lat;
	:northernmost_latitude = +lat;
	:westernmost_longitude = +lon;
	:easternmost_longitude = +lon;
	:quality_statement = "+qual";

data:
    time =  +time;
    latitude = +lat;
    longitude = +lon;
    pres = +pres;
    temp = +temp;
    psal = +psal;
    o2 = +oxygen;
}
