netcdf template_mooring {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 

dimensions:
    time = unlimited;
    n_levels = +nlevels; // maximum number of levels (depth)

variables:
    double time(time);
	time:long_name = "time" ;
	time:short_name = "time" ;
	time:standard_name = "time" ;
	time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
    float depth(n_levels);
	depth:long_name = "Depth in meters";
	depth:short_name = "depth";
	depth:standard_name = "depth";
	depth:units = "meter";
	depth:valid_min = 0;
	depth:valid_max = 15000;
    float latitude;
	latitude:long_name = "latitude";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.f;
	latitude:valid_max = 90.f;
    float longitude;
	longitude:long_name = "longitude";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.f;
	longitude:valid_max = 180.f;
    float pres(time,n_levels);
	pres:long_name = "Sea Water Pressure";
	pres:short_name = "Pressure";
	pres:standard_name = "sea_water_pressure";
	pres:units = "dbar";
	pres:valid_min = 0;
	pres:valid_max = 15000;
    float speed(time,n_levels);
	speed:long_name = "Sea Water Speed";
	speed:short_name = "speed";
	speed:standard_name = "sea_water_speed";
	speed:units = "m s-1";
	speed:valid_min = 0;
	speed:valid_max = 15000;
    float direction(time,n_levels);
	direction:long_name = "Direction of current";
	direction:short_name = "direction";
	direction:standard_name = "direction_of_sea_water_velocity";
	direction:units = "degree";
	direction:valid_min = 0;
	direction:valid_max = 360;
    float ucomp(time,n_levels);
	ucomp:long_name = "Eastwards velocity component of water";
	ucomp:short_name = "eastwards_veolcity";
	ucomp:standard_name = "eastward_sea_water_velocity";
	ucomp:units = "m s-1";
	ucomp:valid_min = 0;
	ucomp:valid_max = 15000;
    float vcomp(time,n_levels);
	vcomp:long_name = "Northwards velocity component of water";
	vcomp:short_name = "northwards_velocity";
	vcomp:standard_name = "northward_sea_water_velocity";
	vcomp:units = "m s-1";
	vcomp:valid_min = 0;
	vcomp:valid_max = 15000;
    float temp(time,n_levels);
	temp:long_name = "Ocean temperature (ITS-90 deg. C)";
	temp:short_name = "temperature";
	temp:_FillValue = 9999.f;
	temp:units = "degrees Celsius";
	temp:valid_min = -3;
	temp:valid_max = 40;
    float psal(time,n_levels);
	psal:long_name = "Practical salinity (PSU/sal00)";
	psal:short_name = "salinity";
	psal:standard_name = "sea_water_salinity";
	psal:_FillValue = 9999.f;
	psal:units = "";
	psal:valid_min = 0;
	psal:valid_max = 60;

// global attributes
	:Conventions = "CF-1.0";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; // Add text if wanted
	:topicCategory = "+topic"; // Blank separated list
	:keywords = "+keyw"; // Blank separated list
	:Area = "+area"; // Comma separated list, see http://damocles.met.no/
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:Product_name = "+pname";
	:Platform_name = "+vessel";
	:start_date = "+start_date";
	:stop_date = "+stop_date";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +lat;
	:northernmost_latitude = +lat;
	:westernmost_longitude = +lon;
	:easternmost_longitude = +lon;

data:
    time =  +time;
    depth = +depth;
    latitude = +lat;
    longitude = +lon;
    pres = +pres;
    speed = +speed;
    direction = +direction;
    ucomp = +ucomp;
    vcomp = +vcomp;
    temp = +temp;
    psal = +psal;
}
