netcdf template_ctd_ugot {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 
// $Id: template_ctd_ugot.cdl,v 1.3 2010-06-16 18:39:52 steingod Exp $
// This template is dedicated for the ISSS08 data delivered by UGOT, it
// basically contains temperature, salinity (and turbidity) at pressure
// levels accompanied by quality flags for each variable and bottom depth
// at the station.

dimensions:
    time = unlimited; //
    n_levels = +ndepths; // maximum number of levels (depth)
    stations = +nstations;
    str25 = 25;

variables:
    char stid(stations,str25);
    	stid:long_name = "Station identifier";
    double time(time);
	time:long_name = "time" ;
	time:short_name = "time" ;
	time:standard_name = "time" ;
	time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
	time:axis = "T";
    float latitude(stations);
	latitude:long_name = "latitude";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.;
	latitude:valid_max = 90.;
    float longitude(stations);
	longitude:long_name = "longitude";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.;
	longitude:valid_max = 180.;
    float bdepth(stations);
	bdepth:long_name = "Depth to ocean bottom";
	bdepth:short_name = "bdepth";
	bdepth:units = "m";
	bdepth:valid_min = 0.;
	bdepth:valid_max = 3000.;
	bdepth:_FillValue = 9999.f;
    float pres(n_levels);
	pres:long_name = "Sea Water Pressure";
	pres:short_name = "Pressure";
	pres:standard_name = "sea_water_pressure";
	pres:units = "dbar";
	pres:valid_min = 0.;
	pres:valid_max = 5000.;
	pres:_FillValue = 9999.f;
	pres:axis = "Y";
    float temp(stations,n_levels);
	temp:long_name = "Ocean temperature (ITS-90 deg. C)";
	temp:short_name = "temperature";
	temp:standard_name = "sea_water_temperature";
	temp:_FillValue = 9999.f;
	temp:units = "degrees Celsius";
	temp:coordinates = "time pres";
	temp:axis = "X";
    float temp_qf(stations,n_levels);
	temp_qf:long_name = "Ocean temperature quality flag (0=OK)";
	temp_qf:short_name = "temperature quality flag";
	temp_qf:_FillValue = 9999.f;
	temp_qf:units = "";
	temp_qf:coordinates = "time pres";
	temp_qf:axis = "X";
    float turb(stations,n_levels);
	turb:long_name = "WET-Labs_ECO_NTU/Turbidity sensor output [V]";
	turb:short_name = "turb";
	turb:_FillValue = 9999.f;
	turb:units = "Volt";
	turb:coordinates = "time pres";
	turb:axis = "X";
    float turb_qf(stations,n_levels);
	turb_qf:long_name = "Ocean turbidity quality flag (0=OK)";
	turb_qf:short_name = "turbidity quality flag";
	turb_qf:_FillValue = 9999.f;
	turb_qf:units = "";
	turb_qf:coordinates = "time pres";
	turb_qf:axis = "X";
    float psal(stations,n_levels);
	psal:long_name = "Practical salinity (PSU/sal00)";
	psal:short_name = "salinity";
	psal:standard_name = "sea_water_salinity";
	psal:_FillValue = 9999.f;
	psal:units = "";
	psal:coordinates = "time pres";
	psal:axis = "X";
    float psal_qf(stations,n_levels);
	psal_qf:long_name = "Ocean salinity quality flag (0=OK)";
	psal_qf:short_name = "salinity quality flag";
	psal_qf:_FillValue = 9999.f;
	psal_qf:units = "";
	psal_qf:coordinates = "time pres";
	psal_qf:axis = "X";

// global attributes
	:Conventions = "CF-1.0";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; // Add text if wanted
	:topiccategory = "+topic"; // Blank separated list
	:keywords = "+keyw"; // Blank separated list
	:gcmd_keywords = "+gcmdkeyw"; // Newline separated list
	:area = "+area"; // Comma separated list, see http://damocles.met.no/
	:activity_type = "+activity";
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:product_name = "+pname";
	:Platform_name = "+vessel";
	:project_name = "+project_name";
	:start_date = "+start_date";
	:stop_date = "+stop_date";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +slat;
	:northernmost_latitude = +nlat;
	:westernmost_longitude = +wlon;
	:easternmost_longitude = +elon;
	:quality_statement = "+qual";
	:operational_status = "+opstatus";

data:
    stid = +stid;
    time =  +time;
    latitude = +lat;
    longitude = +lon;
    bdepth = +bdepth;
    pres = +pres;
    temp = +temp;
    temp_qf = +temp_qf;
    turb = +turb;
    turb_qf = +turb_qf;
    psal = +psal;
    psal_qf = +psal_qf;
}
