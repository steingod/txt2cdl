netcdf template_bio {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 
// $Id: template_seaicethickness.cdl,v 1.1 2011-01-18 14:37:00 steingod Exp $

dimensions:
    time = unlimited;
    stations = +nstations;
    str25 = 25;

variables:
    char stid(stations,str25);
    	stid:long_name = "Station_identifier";
    double time(stations);
	time:long_name = "time_in_UTC_the_station_was_taken";
	time:short_name = "time";
	time:standard_name = "time";
	time:units = "seconds since 1970-01-01 00:00:00 UTC";
	time:axis = "T";
    float latitude(stations);
	latitude:long_name = "geographical_latitude_in_degrees_North";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.;
	latitude:valid_max = 90.;
    float longitude(stations);
	longitude:long_name = "geographical_longitude_in_degrees_East";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.;
	longitude:valid_max = 180.;
    float icet(time);
	icet:standard_name = "sea_ice_thickness";
	icet:long_name = "sea_ice_thickness_in_meter";
	icet:short_name = "icet";
	icet:_FillValue = 9999.f;
	icet:units = "meter";
	icet:coordinates = "time longitude latitude";

// global attributes
	:Conventions = "CF-1.4";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; 
	:topiccategory = "+topic"; 
	:keywords = "+keyw"; 
	:gcmd_keywords = "+gcmdkeyw"; 
	:area = "+area"; 
	:activity_type = "+activity";
	:operational_status = "+opstatus";
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:product_name = "+pname";
	:Platform_name = "+vessel";
	:project_name = "+project_name";
	:start_date = "+start_date";
	:stop_date = "+stop_date";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +slat;
	:northernmost_latitude = +nlat;
	:westernmost_longitude = +wlon;
	:easternmost_longitude = +elon;
	:quality_statement = "+qual";

data:
    stid = +stid;
    time =  +time;
    latitude = +lat;
    longitude = +lon;
    intdepth = +depth;
    icet = +icethickness;
}
