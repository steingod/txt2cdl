netcdf template_itp {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 
// $Id: template_itp.cdl,v 1.1 2008-10-18 21:26:50 steingod Exp $

dimensions:
    time = UNLIMITED; //
    n_levels = +nvalues; // maximum number of levels (depth)

variables:
    double time(time);
	time:long_name = "time" ;
	time:short_name = "time" ;
	time:standard_name = "time" ;
	time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
    float latitude;
	latitude:long_name = "latitude";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.;
	latitude:valid_max = 90.;
    float longitude;
	longitude:long_name = "longitude";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.;
	longitude:valid_max = 180.;
    float pres(n_levels);
	pres:long_name = "Sea Water Pressure";
	pres:short_name = "Pressure";
	pres:standard_name = "sea_water_pressure";
	pres:units = "dbar";
	pres:valid_min = 0.;
	pres:valid_max = 15000.;
    float temp(n_levels);
	temp:long_name = "Ocean temperature (ITS-90 deg. C)";
	temp:short_name = "temperature";
	temp:_FillValue = 9999.f;
	temp:units = "degrees Celsius";
//    char qc_temp(n_levels);
//	qc_temp:long_name = "Quality flag temperature";
//	qc_temp:short_name = "qflgtemp";
//	qc_temp:_FillValue = " ";
    float cond(n_levels);
	cond:long_name = "Ocean conductivity (S/m)";
	cond:short_name = "conductivity";
	cond:standard_name = "sea_water_electrical_conductivity";
	cond:_FillValue = 9999.f;
	cond:units = "S/m";
//    char qc_cond(n_levels);
//	qc_cond:long_name = "Quality flag conductivity";
//	qc_cond:short_name = "qflgcond";
//	qc_cond:_FillValue = " ";
    float psal(n_levels);
	psal:long_name = "Practical salinity (PSU/sal00)";
	psal:short_name = "salinity";
	psal:standard_name = "sea_water_salinity";
	psal:_FillValue = 9999.f;
	psal:units = "";
//    char qc_psal(n_levels);
//	qc_psal:long_name = "Quality flag salinity";
//	qc_psal:short_name = "qflgsal";
//	qc_psal:_FillValue = " ";

// global attributes
	:Conventions = "CF-1.0";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; // Add text if wanted
	:topicCategory = "+topic"; // Blank separated list
	:keywords = "+keyw"; // Blank separated list
	:gcmd_keywords = "+keyw"; // Newline separated list
	:Area = "+area"; // Comma separated list, see http://damocles.met.no/
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:Product_name = "+pname";
	:Platform_name = "+vessel";
	:start_date = "+YYYY-MM-DD HH:MM:SS UTC";
	:stop_date = "+YYYY-MM-DD HH:MM:SS UTC";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +lat;
	:northernmost_latitude = +lat;
	:westernmost_longitude = +lon;
	:easternmost_longitude = +lon;
	:quality_statement = "+qual";

data:
    time =  +time;
    latitude = +lat;
    longitude = +lon;
    pres = +pres;
    temp = +temp;
    cond = +cond;
    psal = +psal;
}
