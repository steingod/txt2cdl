netcdf template_biosediment {

// Template created by �ystein God�y, METNO/FOU, 07.05.2007 
// $Id: template_biosediment.cdl,v 1.4 2010-06-04 12:23:15 steingod Exp $

dimensions:
    depth = +ndepths; 
    stations = +nstations;

variables:
    double time(stations);
	time:long_name = "time in UTC the station was taken";
	time:short_name = "time";
	time:standard_name = "time";
	time:units = "seconds since 1970-01-01 00:00:00 UTC";
	time:axis = "T";
    float latitude(stations);
	latitude:long_name = "geographical latitude in degrees North";
	latitude:short_name = "latitude";
	latitude:standard_name = "latitude";
	latitude:units = "degree_north";
	latitude:valid_min = -90.;
	latitude:valid_max = 90.;
    float longitude(stations);
	longitude:long_name = "geographical longitude in degrees East";
	longitude:short_name = "longitude";
	longitude:standard_name = "longitude";
	longitude:units = "degree_east";
	longitude:valid_min = -180.;
	longitude:valid_max = 180.;
    float depth(depth);
	depth:long_name = "Depth below sea surface in meter";
	depth:short_name = "depth";
	depth:standard_name = "depth";
	depth:units = "m";
	depth:valid_min = 0.;
	depth:valid_max = 15000.;
	depth:positive = "down";
    float chl-a(stations,depth);
	chl-a:long_name = "Chlorophyll-A";
	chl-a:short_name = "chl-a";
	chl-a:_FillValue = 9999.f;
	chl-a:units = "milligram m-2 day-1";
	chl-a:coordinates = "time longitude latitude depth";
    float chl-a_stdev(stations,depth);
	chl-a_stdev:long_name = "Chlorophyll-A standard deviation";
	chl-a_stdev:short_name = "chl-a stdev";
	chl-a_stdev:_FillValue = 9999.f;
	chl-a_stdev:units = "milligram m-2 day-2";
	chl-a_stdev:coordinates = "time longitude latitude depth";
    float phaeopigment(stations,depth);
	phaeopigment:long_name = "Phaeopigment";
	phaeopigment:short_name = "phaeopigment";
	phaeopigment:_FillValue = 9999.f;
	phaeopigment:units = "milligram m-2 day-1";
	phaeopigment:coordinates = "time longitude latitude depth";
    float phaeopigment_stdev(stations,depth);
	phaeopigment_stdev:long_name = "Phaeopigment standard deviation";
	phaeopigment_stdev:short_name = "phaeopigment stdev";
	phaeopigment_stdev:_FillValue = 9999.f;
	phaeopigment_stdev:units = "milligram m-2 day-1";
	phaeopigment_stdev:coordinates = "time longitude latitude depth";
    float POC(stations,depth);
	POC:long_name = "Particulate Organic Carbon";
	POC:short_name = "POC";
	POC:_FillValue = 9999.f;
	POC:units = "milligram m-2 day-1";
	POC:coordinates = "time longitude latitude depth";
    float POC_stdev(stations,depth);
	POC_stdev:long_name = "Particulate Organic Carbon standard deviation";
	POC_stdev:short_name = "POC_stdev";
	POC_stdev:_FillValue = 9999.f;
	POC_stdev:units = "milligram m-2 day-1";
	POC_stdev:coordinates = "time longitude latitude depth";
    float PON(stations,depth);
	PON:long_name = "Particulate Organic Nitrogen";
	PON:short_name = "PON";
	PON:_FillValue = 9999.f;
	PON:units = "milligram m-2 day-1";
	PON:coordinates = "time longitude latitude depth";
    float PON_stdev(stations,depth);
	PON_stdev:long_name = "Particulate Organic Nitrogen standard deviation";
	PON_stdev:short_name = "PON_stdev";
	PON_stdev:_FillValue = 9999.f;
	PON_stdev:units = "milligram m-2 day-1";
	PON_stdev:coordinates = "time longitude latitude depth";
    float FPC(stations,depth);
	FPC:long_name = "Feacal Pellet Carbon";
	FPC:short_name = "FPC";
	FPC:_FillValue = 9999.f;
	FPC:units = "milligram m-2 day-1";
	FPC:coordinates = "time longitude latitude depth";

// global attributes
	:Conventions = "CF-1.4";
	:history = "+history";
	:title = "+title";
	:abstract = "+abstract"; 
	:topiccategory = "+topic"; 
	:keywords = "+keyw"; 
	:gcmd_keywords = "+gcmdkeyw"; 
	:area = "+area"; 
	:activity_type = "+activity";
	:operational_status = "+opstatus";
	:PI_name = "+piname";
	:contact = "+email";
	:institution = "+inst";
	:url = "+url";
	:product_name = "+pname";
	:Platform_name = "+vessel";
	:project_name = "+project_name";
	:start_date = "+start_date";
	:stop_date = "+stop_date";
	:distribution_statement = "+distribution"; 
	:southernmost_latitude = +slat;
	:northernmost_latitude = +nlat;
	:westernmost_longitude = +wlon;
	:easternmost_longitude = +elon;
	:quality_statement = "+qual";

data:
    time =  +time;
    latitude = +lat;
    longitude = +lon;
    depth = +depth;
    chl-a = +chl-a;
    chl-a_stdev = +chl-a_stdev;
    phaeopigment = +pigm;
    phaeopigment_stdev = +pigm_stdev;
    POC = +poc;
    POC_stdev = +poc_stdev;
    PON = +pon;
    PON_stdev = +pon_stdev;
    FPC = +fpc;
}
